//FC0_node0
wire signed[15:0] fc0_node0_c[29:0];
assign fc0_node0_c[0] = 16'h0292;
assign fc0_node0_c[1] = 16'h0091;
assign fc0_node0_c[2] = 16'hFD77;
assign fc0_node0_c[3] = 16'h0045;
assign fc0_node0_c[4] = 16'hFE45;
assign fc0_node0_c[5] = 16'hFD24;
assign fc0_node0_c[6] = 16'h0297;
assign fc0_node0_c[7] = 16'h0238;
assign fc0_node0_c[8] = 16'hFD18;
assign fc0_node0_c[9] = 16'h008C;
assign fc0_node0_c[10] = 16'hFF82;
assign fc0_node0_c[11] = 16'hFF86;
assign fc0_node0_c[12] = 16'hFEAD;
assign fc0_node0_c[13] = 16'h0128;
assign fc0_node0_c[14] = 16'hFE48;
assign fc0_node0_c[15] = 16'h0A31;
assign fc0_node0_c[16] = 16'h0520;
assign fc0_node0_c[17] = 16'hFE27;
assign fc0_node0_c[18] = 16'hFCED;
assign fc0_node0_c[19] = 16'hFDF6;
assign fc0_node0_c[20] = 16'hF821;
assign fc0_node0_c[21] = 16'hFE4B;
assign fc0_node0_c[22] = 16'hFDA0;
assign fc0_node0_c[23] = 16'h01BE;
assign fc0_node0_c[24] = 16'h054E;
assign fc0_node0_c[25] = 16'h02F9;
assign fc0_node0_c[26] = 16'h05BB;
assign fc0_node0_c[27] = 16'h0329;
assign fc0_node0_c[28] = 16'h0320;
assign fc0_node0_c[29] = 16'h0142;


//FC0_node1
wire signed[15:0] fc0_node1_c[29:0];
assign fc0_node1_c[0] = 16'hFFF3;
assign fc0_node1_c[1] = 16'hFDCC;
assign fc0_node1_c[2] = 16'hFDC0;
assign fc0_node1_c[3] = 16'hFFD8;
assign fc0_node1_c[4] = 16'h0074;
assign fc0_node1_c[5] = 16'hFEAF;
assign fc0_node1_c[6] = 16'h01BB;
assign fc0_node1_c[7] = 16'hFE3B;
assign fc0_node1_c[8] = 16'h02A5;
assign fc0_node1_c[9] = 16'h0200;
assign fc0_node1_c[10] = 16'hFD8B;
assign fc0_node1_c[11] = 16'hFF47;
assign fc0_node1_c[12] = 16'h0022;
assign fc0_node1_c[13] = 16'h0072;
assign fc0_node1_c[14] = 16'h00B2;
assign fc0_node1_c[15] = 16'h176F;
assign fc0_node1_c[16] = 16'h07DB;
assign fc0_node1_c[17] = 16'hF423;
assign fc0_node1_c[18] = 16'h049B;
assign fc0_node1_c[19] = 16'hF8ED;
assign fc0_node1_c[20] = 16'hF61D;
assign fc0_node1_c[21] = 16'hFBDC;
assign fc0_node1_c[22] = 16'hF95F;
assign fc0_node1_c[23] = 16'h009C;
assign fc0_node1_c[24] = 16'h02ED;
assign fc0_node1_c[25] = 16'hFE48;
assign fc0_node1_c[26] = 16'h03C2;
assign fc0_node1_c[27] = 16'h0026;
assign fc0_node1_c[28] = 16'hFFE5;
assign fc0_node1_c[29] = 16'h00E8;


//FC0_node2
wire signed[15:0] fc0_node2_c[29:0];
assign fc0_node2_c[0] = 16'hFFB4;
assign fc0_node2_c[1] = 16'h0011;
assign fc0_node2_c[2] = 16'hFFC0;
assign fc0_node2_c[3] = 16'h0097;
assign fc0_node2_c[4] = 16'h01DB;
assign fc0_node2_c[5] = 16'h0295;
assign fc0_node2_c[6] = 16'h01DA;
assign fc0_node2_c[7] = 16'h02C6;
assign fc0_node2_c[8] = 16'hFFCB;
assign fc0_node2_c[9] = 16'hFD62;
assign fc0_node2_c[10] = 16'hFE9F;
assign fc0_node2_c[11] = 16'h01FC;
assign fc0_node2_c[12] = 16'hFFFD;
assign fc0_node2_c[13] = 16'hFE8B;
assign fc0_node2_c[14] = 16'hFDC4;
assign fc0_node2_c[15] = 16'h0478;
assign fc0_node2_c[16] = 16'h0320;
assign fc0_node2_c[17] = 16'h0456;
assign fc0_node2_c[18] = 16'hECD0;
assign fc0_node2_c[19] = 16'h0CD5;
assign fc0_node2_c[20] = 16'h0024;
assign fc0_node2_c[21] = 16'hF2D8;
assign fc0_node2_c[22] = 16'h05CB;
assign fc0_node2_c[23] = 16'h09DF;
assign fc0_node2_c[24] = 16'h1222;
assign fc0_node2_c[25] = 16'hFE3C;
assign fc0_node2_c[26] = 16'h0082;
assign fc0_node2_c[27] = 16'hFA7B;
assign fc0_node2_c[28] = 16'hFF83;
assign fc0_node2_c[29] = 16'h0741;


//FC0_node3
wire signed[15:0] fc0_node3_c[29:0];
assign fc0_node3_c[0] = 16'h0009;
assign fc0_node3_c[1] = 16'hFEAB;
assign fc0_node3_c[2] = 16'h0119;
assign fc0_node3_c[3] = 16'hFD60;
assign fc0_node3_c[4] = 16'hFFBB;
assign fc0_node3_c[5] = 16'h0278;
assign fc0_node3_c[6] = 16'hFED0;
assign fc0_node3_c[7] = 16'h02A2;
assign fc0_node3_c[8] = 16'h010D;
assign fc0_node3_c[9] = 16'hFD5E;
assign fc0_node3_c[10] = 16'h01D8;
assign fc0_node3_c[11] = 16'hFFAA;
assign fc0_node3_c[12] = 16'hFEB2;
assign fc0_node3_c[13] = 16'h0250;
assign fc0_node3_c[14] = 16'hFDA3;
assign fc0_node3_c[15] = 16'hFD96;
assign fc0_node3_c[16] = 16'h01CC;
assign fc0_node3_c[17] = 16'h0B56;
assign fc0_node3_c[18] = 16'hE647;
assign fc0_node3_c[19] = 16'h0F83;
assign fc0_node3_c[20] = 16'h0EE8;
assign fc0_node3_c[21] = 16'hFB97;
assign fc0_node3_c[22] = 16'h04DB;
assign fc0_node3_c[23] = 16'h03C6;
assign fc0_node3_c[24] = 16'h05A4;
assign fc0_node3_c[25] = 16'h015F;
assign fc0_node3_c[26] = 16'h084E;
assign fc0_node3_c[27] = 16'h0866;
assign fc0_node3_c[28] = 16'hFF6B;
assign fc0_node3_c[29] = 16'h01AD;


//FC0_node4
wire signed[15:0] fc0_node4_c[29:0];
assign fc0_node4_c[0] = 16'hFE66;
assign fc0_node4_c[1] = 16'hFE50;
assign fc0_node4_c[2] = 16'h00FF;
assign fc0_node4_c[3] = 16'hFE43;
assign fc0_node4_c[4] = 16'hFFE4;
assign fc0_node4_c[5] = 16'h0038;
assign fc0_node4_c[6] = 16'h01E1;
assign fc0_node4_c[7] = 16'hFDCD;
assign fc0_node4_c[8] = 16'hFE02;
assign fc0_node4_c[9] = 16'hFE4F;
assign fc0_node4_c[10] = 16'h020B;
assign fc0_node4_c[11] = 16'hFEF4;
assign fc0_node4_c[12] = 16'h0274;
assign fc0_node4_c[13] = 16'h0108;
assign fc0_node4_c[14] = 16'h005E;
assign fc0_node4_c[15] = 16'hF0C5;
assign fc0_node4_c[16] = 16'h007A;
assign fc0_node4_c[17] = 16'h0AF5;
assign fc0_node4_c[18] = 16'h04DF;
assign fc0_node4_c[19] = 16'hFD4E;
assign fc0_node4_c[20] = 16'hEFB7;
assign fc0_node4_c[21] = 16'h016E;
assign fc0_node4_c[22] = 16'hFEF5;
assign fc0_node4_c[23] = 16'h0397;
assign fc0_node4_c[24] = 16'h0836;
assign fc0_node4_c[25] = 16'h0932;
assign fc0_node4_c[26] = 16'h08D3;
assign fc0_node4_c[27] = 16'hFCE7;
assign fc0_node4_c[28] = 16'hFF8A;
assign fc0_node4_c[29] = 16'h0233;


//FC0_node5
wire signed[15:0] fc0_node5_c[29:0];
assign fc0_node5_c[0] = 16'h0172;
assign fc0_node5_c[1] = 16'hFDEF;
assign fc0_node5_c[2] = 16'hFF2C;
assign fc0_node5_c[3] = 16'hFF05;
assign fc0_node5_c[4] = 16'hFF7E;
assign fc0_node5_c[5] = 16'h0021;
assign fc0_node5_c[6] = 16'h0268;
assign fc0_node5_c[7] = 16'h005D;
assign fc0_node5_c[8] = 16'h029D;
assign fc0_node5_c[9] = 16'h01C8;
assign fc0_node5_c[10] = 16'hFE28;
assign fc0_node5_c[11] = 16'h014F;
assign fc0_node5_c[12] = 16'hFDEE;
assign fc0_node5_c[13] = 16'hFEC0;
assign fc0_node5_c[14] = 16'h00DA;
assign fc0_node5_c[15] = 16'hF6AC;
assign fc0_node5_c[16] = 16'h04F9;
assign fc0_node5_c[17] = 16'h0634;
assign fc0_node5_c[18] = 16'h024A;
assign fc0_node5_c[19] = 16'h0020;
assign fc0_node5_c[20] = 16'hF202;
assign fc0_node5_c[21] = 16'h0E8A;
assign fc0_node5_c[22] = 16'hF823;
assign fc0_node5_c[23] = 16'hFE7D;
assign fc0_node5_c[24] = 16'hFEFC;
assign fc0_node5_c[25] = 16'h0833;
assign fc0_node5_c[26] = 16'h0E80;
assign fc0_node5_c[27] = 16'h0D53;
assign fc0_node5_c[28] = 16'hFEE1;
assign fc0_node5_c[29] = 16'h0085;


//FC0_node6
wire signed[15:0] fc0_node6_c[29:0];
assign fc0_node6_c[0] = 16'hFEED;
assign fc0_node6_c[1] = 16'hFD1E;
assign fc0_node6_c[2] = 16'h0151;
assign fc0_node6_c[3] = 16'hFE99;
assign fc0_node6_c[4] = 16'hFE17;
assign fc0_node6_c[5] = 16'hFE63;
assign fc0_node6_c[6] = 16'h01AD;
assign fc0_node6_c[7] = 16'h018C;
assign fc0_node6_c[8] = 16'h023F;
assign fc0_node6_c[9] = 16'h010F;
assign fc0_node6_c[10] = 16'hFF07;
assign fc0_node6_c[11] = 16'hFF30;
assign fc0_node6_c[12] = 16'h00DC;
assign fc0_node6_c[13] = 16'h0264;
assign fc0_node6_c[14] = 16'h00CC;
assign fc0_node6_c[15] = 16'hFD32;
assign fc0_node6_c[16] = 16'hFE73;
assign fc0_node6_c[17] = 16'hFB27;
assign fc0_node6_c[18] = 16'h161D;
assign fc0_node6_c[19] = 16'hF7DA;
assign fc0_node6_c[20] = 16'hED75;
assign fc0_node6_c[21] = 16'h0059;
assign fc0_node6_c[22] = 16'hFCA8;
assign fc0_node6_c[23] = 16'hFAC6;
assign fc0_node6_c[24] = 16'h0622;
assign fc0_node6_c[25] = 16'h037B;
assign fc0_node6_c[26] = 16'hF778;
assign fc0_node6_c[27] = 16'hED7D;
assign fc0_node6_c[28] = 16'h01D5;
assign fc0_node6_c[29] = 16'h005A;


//FC0_node7
wire signed[15:0] fc0_node7_c[29:0];
assign fc0_node7_c[0] = 16'h026C;
assign fc0_node7_c[1] = 16'hFF0A;
assign fc0_node7_c[2] = 16'h00DC;
assign fc0_node7_c[3] = 16'hFF55;
assign fc0_node7_c[4] = 16'hFFE4;
assign fc0_node7_c[5] = 16'hFE63;
assign fc0_node7_c[6] = 16'h00FC;
assign fc0_node7_c[7] = 16'h00EC;
assign fc0_node7_c[8] = 16'hFFF2;
assign fc0_node7_c[9] = 16'hFF59;
assign fc0_node7_c[10] = 16'hFE34;
assign fc0_node7_c[11] = 16'h0204;
assign fc0_node7_c[12] = 16'hFDD3;
assign fc0_node7_c[13] = 16'h012C;
assign fc0_node7_c[14] = 16'hFF04;
assign fc0_node7_c[15] = 16'hEF44;
assign fc0_node7_c[16] = 16'hFC56;
assign fc0_node7_c[17] = 16'h053C;
assign fc0_node7_c[18] = 16'h0603;
assign fc0_node7_c[19] = 16'h01DD;
assign fc0_node7_c[20] = 16'hFCD1;
assign fc0_node7_c[21] = 16'h024F;
assign fc0_node7_c[22] = 16'h049C;
assign fc0_node7_c[23] = 16'hFFE4;
assign fc0_node7_c[24] = 16'h0145;
assign fc0_node7_c[25] = 16'h0169;
assign fc0_node7_c[26] = 16'hFC6C;
assign fc0_node7_c[27] = 16'hF99F;
assign fc0_node7_c[28] = 16'hFF3F;
assign fc0_node7_c[29] = 16'h02EA;


//FC0_node8
wire signed[15:0] fc0_node8_c[29:0];
assign fc0_node8_c[0] = 16'h01F2;
assign fc0_node8_c[1] = 16'hFE7C;
assign fc0_node8_c[2] = 16'h0007;
assign fc0_node8_c[3] = 16'h0135;
assign fc0_node8_c[4] = 16'h0041;
assign fc0_node8_c[5] = 16'h0057;
assign fc0_node8_c[6] = 16'h005D;
assign fc0_node8_c[7] = 16'hFDB5;
assign fc0_node8_c[8] = 16'h003B;
assign fc0_node8_c[9] = 16'h0205;
assign fc0_node8_c[10] = 16'h02A1;
assign fc0_node8_c[11] = 16'h01B7;
assign fc0_node8_c[12] = 16'h0063;
assign fc0_node8_c[13] = 16'h0152;
assign fc0_node8_c[14] = 16'hFE94;
assign fc0_node8_c[15] = 16'hE176;
assign fc0_node8_c[16] = 16'hF481;
assign fc0_node8_c[17] = 16'h1015;
assign fc0_node8_c[18] = 16'h0402;
assign fc0_node8_c[19] = 16'h0801;
assign fc0_node8_c[20] = 16'h053D;
assign fc0_node8_c[21] = 16'hFF1A;
assign fc0_node8_c[22] = 16'h0A0A;
assign fc0_node8_c[23] = 16'hFE93;
assign fc0_node8_c[24] = 16'h0288;
assign fc0_node8_c[25] = 16'h01A5;
assign fc0_node8_c[26] = 16'hF6B2;
assign fc0_node8_c[27] = 16'hF50B;
assign fc0_node8_c[28] = 16'h01A3;
assign fc0_node8_c[29] = 16'h0139;


//FC1_node0
wire signed[15:0] fc1_node0_c[8:0];
assign fc1_node0_c[0] = 16'hFFEC;
assign fc1_node0_c[1] = 16'h092C;
assign fc1_node0_c[2] = 16'hFC3E;
assign fc1_node0_c[3] = 16'hEA17;
assign fc1_node0_c[4] = 16'h0404;
assign fc1_node0_c[5] = 16'hF80F;
assign fc1_node0_c[6] = 16'h1BAB;
assign fc1_node0_c[7] = 16'h0380;
assign fc1_node0_c[8] = 16'h0550;


//FC1_node1
wire signed[15:0] fc1_node1_c[8:0];
assign fc1_node1_c[0] = 16'h035F;
assign fc1_node1_c[1] = 16'h0A78;
assign fc1_node1_c[2] = 16'hED79;
assign fc1_node1_c[3] = 16'hF59A;
assign fc1_node1_c[4] = 16'hFB2E;
assign fc1_node1_c[5] = 16'h0B31;
assign fc1_node1_c[6] = 16'h00D0;
assign fc1_node1_c[7] = 16'hF7C5;
assign fc1_node1_c[8] = 16'hF0A5;


//FC1_node2
wire signed[15:0] fc1_node2_c[8:0];
assign fc1_node2_c[0] = 16'hFB2A;
assign fc1_node2_c[1] = 16'hFA58;
assign fc1_node2_c[2] = 16'h0AE2;
assign fc1_node2_c[3] = 16'h0EE8;
assign fc1_node2_c[4] = 16'hF292;
assign fc1_node2_c[5] = 16'hEFA9;
assign fc1_node2_c[6] = 16'hF48F;
assign fc1_node2_c[7] = 16'hFC4B;
assign fc1_node2_c[8] = 16'h0802;


//FC1_node3
wire signed[15:0] fc1_node3_c[8:0];
assign fc1_node3_c[0] = 16'hFADC;
assign fc1_node3_c[1] = 16'hEEB3;
assign fc1_node3_c[2] = 16'hFBEB;
assign fc1_node3_c[3] = 16'h07D4;
assign fc1_node3_c[4] = 16'h0A79;
assign fc1_node3_c[5] = 16'h0BFA;
assign fc1_node3_c[6] = 16'hFC1F;
assign fc1_node3_c[7] = 16'h0895;
assign fc1_node3_c[8] = 16'h161C;


//FC1_node4
wire signed[15:0] fc1_node4_c[8:0];
assign fc1_node4_c[0] = 16'h0B3E;
assign fc1_node4_c[1] = 16'h0AC8;
assign fc1_node4_c[2] = 16'h152E;
assign fc1_node4_c[3] = 16'h0BD6;
assign fc1_node4_c[4] = 16'h0684;
assign fc1_node4_c[5] = 16'h03F1;
assign fc1_node4_c[6] = 16'hF9AB;
assign fc1_node4_c[7] = 16'hF86F;
assign fc1_node4_c[8] = 16'hF4B6;


