reg [31:0] FIR_C0 = 32'h0000B203;    // 0.00016976520419120789
reg [31:0] FIR_C1 = 32'h00003181;    // 0.00004721060395240784
reg [31:0] FIR_C2 = 32'hFFFF864B;    // -0.00011606886982917786
reg [31:0] FIR_C3 = 32'hFFFED465;    // -0.00028572604060173035
reg [31:0] FIR_C4 = 32'hFFFEE129;    // -0.00027355179190635681
reg [31:0] FIR_C5 = 32'h000008F9;    // 0.00000855699181556702
reg [31:0] FIR_C6 = 32'h0001A798;    // 0.00040397047996520996
reg [31:0] FIR_C7 = 32'h00024FF6;    // 0.00056453794240951538
reg [31:0] FIR_C8 = 32'h0000F1CA;    // 0.00023058801889419556
reg [31:0] FIR_C9 = 32'hFFFE1436;    // -0.00046900659799575806
reg [31:0] FIR_C10 = 32'hFFFBEE58;    // -0.00099340081214904785
reg [31:0] FIR_C11 = 32'hFFFCD644;    // -0.00077222287654876709
reg [31:0] FIR_C12 = 32'h0001036E;    // 0.00024741142988204956
reg [31:0] FIR_C13 = 32'h00059FCA;    // 0.00137308984994888306
reg [31:0] FIR_C14 = 32'h00067ED1;    // 0.00158578529953956604
reg [31:0] FIR_C15 = 32'h0001A7AB;    // 0.00040404126048088074
reg [31:0] FIR_C16 = 32'hFFF9DBAF;    // -0.00149947777390480042
reg [31:0] FIR_C17 = 32'hFFF566C7;    // -0.00258753076195716858
reg [31:0] FIR_C18 = 32'hFFF949BF;    // -0.00163865461945533752
reg [31:0] FIR_C19 = 32'h000442E3;    // 0.00104035064578056335
reg [31:0] FIR_C20 = 32'h000E4861;    // 0.00348699465394020081
reg [31:0] FIR_C21 = 32'h000E18D4;    // 0.00344164669513702393
reg [31:0] FIR_C22 = 32'h00015094;    // 0.00032098591327667236
reg [31:0] FIR_C23 = 32'hFFF04341;    // -0.00384211167693138123
reg [31:0] FIR_C24 = 32'hFFE91589;    // -0.00559469684958457947
reg [31:0] FIR_C25 = 32'hFFF4752F;    // -0.00281793251633644104
reg [31:0] FIR_C26 = 32'h000C9948;    // 0.00307586789131164551
reg [31:0] FIR_C27 = 32'h001F1C74;    // 0.00759549438953399658
reg [31:0] FIR_C28 = 32'h001A729E;    // 0.00645696371793746948
reg [31:0] FIR_C29 = 32'hFFFD943B;    // -0.00059105828404426575
reg [31:0] FIR_C30 = 32'hFFDC8104;    // -0.00866602361202239990
reg [31:0] FIR_C31 = 32'hFFD342CF;    // -0.01092261448502540588
reg [31:0] FIR_C32 = 32'hFFEF2149;    // -0.00411864742636680603
reg [31:0] FIR_C33 = 32'h001FDF2C;    // 0.00778119266033172607
reg [31:0] FIR_C34 = 32'h003F8169;    // 0.01550427451729774475
reg [31:0] FIR_C35 = 32'h002E9588;    // 0.01137307286262512207
reg [31:0] FIR_C36 = 32'hFFF0DF30;    // -0.00369340181350708008
reg [31:0] FIR_C37 = 32'hFFB1ED1B;    // -0.01906098797917366028
reg [31:0] FIR_C38 = 32'hFFA89835;    // -0.02133921906352043152
reg [31:0] FIR_C39 = 32'hFFEA81BB;    // -0.00524737313389778137
reg [31:0] FIR_C40 = 32'h00517CAA;    // 0.01989427953958511353
reg [31:0] FIR_C41 = 32'h008CEDEC;    // 0.03440658748149871826
reg [31:0] FIR_C42 = 32'h005AB35B;    // 0.02214370295405387878
reg [31:0] FIR_C43 = 32'hFFC2B5A1;    // -0.01496350392699241638
reg [31:0] FIR_C44 = 32'hFF272F92;    // -0.05293314903974533081
reg [31:0] FIR_C45 = 32'hFF147F7A;    // -0.05749561637639999390
reg [31:0] FIR_C46 = 32'hFFE7CF85;    // -0.00590560957789421082
reg [31:0] FIR_C47 = 32'h01853667;    // 0.09502258524298667908
reg [31:0] FIR_C48 = 32'h035259BC;    // 0.20760510861873626709
reg [31:0] FIR_C49 = 32'h04812148;    // 0.28152588009834289551
reg [31:0] FIR_C50 = 32'h04812148;    // 0.28152588009834289551
reg [31:0] FIR_C51 = 32'h035259BC;    // 0.20760510861873626709
reg [31:0] FIR_C52 = 32'h01853667;    // 0.09502258524298667908
reg [31:0] FIR_C53 = 32'hFFE7CF85;    // -0.00590560957789421082
reg [31:0] FIR_C54 = 32'hFF147F7A;    // -0.05749561637639999390
reg [31:0] FIR_C55 = 32'hFF272F92;    // -0.05293314903974533081
reg [31:0] FIR_C56 = 32'hFFC2B5A1;    // -0.01496350392699241638
reg [31:0] FIR_C57 = 32'h005AB35B;    // 0.02214370295405387878
reg [31:0] FIR_C58 = 32'h008CEDEC;    // 0.03440658748149871826
reg [31:0] FIR_C59 = 32'h00517CAA;    // 0.01989427953958511353
reg [31:0] FIR_C60 = 32'hFFEA81BB;    // -0.00524737313389778137
reg [31:0] FIR_C61 = 32'hFFA89835;    // -0.02133921906352043152
reg [31:0] FIR_C62 = 32'hFFB1ED1B;    // -0.01906098797917366028
reg [31:0] FIR_C63 = 32'hFFF0DF30;    // -0.00369340181350708008
reg [31:0] FIR_C64 = 32'h002E9588;    // 0.01137307286262512207
reg [31:0] FIR_C65 = 32'h003F8169;    // 0.01550427451729774475
reg [31:0] FIR_C66 = 32'h001FDF2C;    // 0.00778119266033172607
reg [31:0] FIR_C67 = 32'hFFEF2149;    // -0.00411864742636680603
reg [31:0] FIR_C68 = 32'hFFD342CF;    // -0.01092261448502540588
reg [31:0] FIR_C69 = 32'hFFDC8104;    // -0.00866602361202239990
reg [31:0] FIR_C70 = 32'hFFFD943B;    // -0.00059105828404426575
reg [31:0] FIR_C71 = 32'h001A729E;    // 0.00645696371793746948
reg [31:0] FIR_C72 = 32'h001F1C74;    // 0.00759549438953399658
reg [31:0] FIR_C73 = 32'h000C9948;    // 0.00307586789131164551
reg [31:0] FIR_C74 = 32'hFFF4752F;    // -0.00281793251633644104
reg [31:0] FIR_C75 = 32'hFFE91589;    // -0.00559469684958457947
reg [31:0] FIR_C76 = 32'hFFF04341;    // -0.00384211167693138123
reg [31:0] FIR_C77 = 32'h00015094;    // 0.00032098591327667236
reg [31:0] FIR_C78 = 32'h000E18D4;    // 0.00344164669513702393
reg [31:0] FIR_C79 = 32'h000E4861;    // 0.00348699465394020081
reg [31:0] FIR_C80 = 32'h000442E3;    // 0.00104035064578056335
reg [31:0] FIR_C81 = 32'hFFF949BF;    // -0.00163865461945533752
reg [31:0] FIR_C82 = 32'hFFF566C7;    // -0.00258753076195716858
reg [31:0] FIR_C83 = 32'hFFF9DBAF;    // -0.00149947777390480042
reg [31:0] FIR_C84 = 32'h0001A7AB;    // 0.00040404126048088074
reg [31:0] FIR_C85 = 32'h00067ED1;    // 0.00158578529953956604
reg [31:0] FIR_C86 = 32'h00059FCA;    // 0.00137308984994888306
reg [31:0] FIR_C87 = 32'h0001036E;    // 0.00024741142988204956
reg [31:0] FIR_C88 = 32'hFFFCD644;    // -0.00077222287654876709
reg [31:0] FIR_C89 = 32'hFFFBEE58;    // -0.00099340081214904785
reg [31:0] FIR_C90 = 32'hFFFE1436;    // -0.00046900659799575806
reg [31:0] FIR_C91 = 32'h0000F1CA;    // 0.00023058801889419556
reg [31:0] FIR_C92 = 32'h00024FF6;    // 0.00056453794240951538
reg [31:0] FIR_C93 = 32'h0001A798;    // 0.00040397047996520996
reg [31:0] FIR_C94 = 32'h000008F9;    // 0.00000855699181556702
reg [31:0] FIR_C95 = 32'hFFFEE129;    // -0.00027355179190635681
reg [31:0] FIR_C96 = 32'hFFFED465;    // -0.00028572604060173035
reg [31:0] FIR_C97 = 32'hFFFF864B;    // -0.00011606886982917786
reg [31:0] FIR_C98 = 32'h00003181;    // 0.00004721060395240784
reg [31:0] FIR_C99 = 32'h0000B203;    // 0.00016976520419120789
