//conv0 kernel0 coeff
wire signed[15:0] conv0_kernel0_c[4:0];
assign conv0_kernel0_c[0] = 16'hE8E7;
assign conv0_kernel0_c[1] = 16'hF728;
assign conv0_kernel0_c[2] = 16'hF47A;
assign conv0_kernel0_c[3] = 16'hF677;
assign conv0_kernel0_c[4] = 16'hF8D5;


//conv0 kernel1 coeff
wire signed[15:0] conv0_kernel1_c[4:0];
assign conv0_kernel1_c[0] = 16'h0591;
assign conv0_kernel1_c[1] = 16'h0341;
assign conv0_kernel1_c[2] = 16'h07B8;
assign conv0_kernel1_c[3] = 16'h0938;
assign conv0_kernel1_c[4] = 16'h2832;


//conv0 kernel2 coeff
wire signed[15:0] conv0_kernel2_c[4:0];
assign conv0_kernel2_c[0] = 16'hE5E9;
assign conv0_kernel2_c[1] = 16'hF2E0;
assign conv0_kernel2_c[2] = 16'hF6AF;
assign conv0_kernel2_c[3] = 16'hFC48;
assign conv0_kernel2_c[4] = 16'hFF99;


//conv0 kernel3 coeff
wire signed[15:0] conv0_kernel3_c[4:0];
assign conv0_kernel3_c[0] = 16'hF793;
assign conv0_kernel3_c[1] = 16'hFDE1;
assign conv0_kernel3_c[2] = 16'h01E8;
assign conv0_kernel3_c[3] = 16'hF949;
assign conv0_kernel3_c[4] = 16'hFB15;


//conv0 kernel4 coeff
wire signed[15:0] conv0_kernel4_c[4:0];
assign conv0_kernel4_c[0] = 16'h00A4;
assign conv0_kernel4_c[1] = 16'h0386;
assign conv0_kernel4_c[2] = 16'hFC1B;
assign conv0_kernel4_c[3] = 16'h090C;
assign conv0_kernel4_c[4] = 16'h161A;


//conv1 kernel0_0 coeff
wire signed[15:0] conv1_kernel0_0_c[4:0];
assign conv1_kernel0_0_c[0] = 16'h0054;
assign conv1_kernel0_0_c[1] = 16'h029F;
assign conv1_kernel0_0_c[2] = 16'hFCBF;
assign conv1_kernel0_0_c[3] = 16'hFD7F;
assign conv1_kernel0_0_c[4] = 16'hFEC5;


//conv1 kernel0_1 coeff
wire signed[15:0] conv1_kernel0_1_c[4:0];
assign conv1_kernel0_1_c[0] = 16'hFE55;
assign conv1_kernel0_1_c[1] = 16'h023F;
assign conv1_kernel0_1_c[2] = 16'hFD7B;
assign conv1_kernel0_1_c[3] = 16'hFE79;
assign conv1_kernel0_1_c[4] = 16'hFDC4;


//conv1 kernel0_2 coeff
wire signed[15:0] conv1_kernel0_2_c[4:0];
assign conv1_kernel0_2_c[0] = 16'hFCFE;
assign conv1_kernel0_2_c[1] = 16'hFDD3;
assign conv1_kernel0_2_c[2] = 16'h0241;
assign conv1_kernel0_2_c[3] = 16'h00B8;
assign conv1_kernel0_2_c[4] = 16'h00D1;


//conv1 kernel0_3 coeff
wire signed[15:0] conv1_kernel0_3_c[4:0];
assign conv1_kernel0_3_c[0] = 16'h0017;
assign conv1_kernel0_3_c[1] = 16'hFE39;
assign conv1_kernel0_3_c[2] = 16'h0067;
assign conv1_kernel0_3_c[3] = 16'hFCD9;
assign conv1_kernel0_3_c[4] = 16'hFDA4;


//conv1 kernel0_4 coeff
wire signed[15:0] conv1_kernel0_4_c[4:0];
assign conv1_kernel0_4_c[0] = 16'hFDF4;
assign conv1_kernel0_4_c[1] = 16'h0181;
assign conv1_kernel0_4_c[2] = 16'h016A;
assign conv1_kernel0_4_c[3] = 16'hFE72;
assign conv1_kernel0_4_c[4] = 16'hFFE0;


//conv1 kernel1_0 coeff
wire signed[15:0] conv1_kernel1_0_c[4:0];
assign conv1_kernel1_0_c[0] = 16'hF51F;
assign conv1_kernel1_0_c[1] = 16'h187F;
assign conv1_kernel1_0_c[2] = 16'h0F60;
assign conv1_kernel1_0_c[3] = 16'hFB33;
assign conv1_kernel1_0_c[4] = 16'hF4FA;


//conv1 kernel1_1 coeff
wire signed[15:0] conv1_kernel1_1_c[4:0];
assign conv1_kernel1_1_c[0] = 16'hF3C7;
assign conv1_kernel1_1_c[1] = 16'h097B;
assign conv1_kernel1_1_c[2] = 16'hF0C1;
assign conv1_kernel1_1_c[3] = 16'hDD71;
assign conv1_kernel1_1_c[4] = 16'h2566;


//conv1 kernel1_2 coeff
wire signed[15:0] conv1_kernel1_2_c[4:0];
assign conv1_kernel1_2_c[0] = 16'hEF80;
assign conv1_kernel1_2_c[1] = 16'h18E3;
assign conv1_kernel1_2_c[2] = 16'h0ED7;
assign conv1_kernel1_2_c[3] = 16'h001F;
assign conv1_kernel1_2_c[4] = 16'hF521;


//conv1 kernel1_3 coeff
wire signed[15:0] conv1_kernel1_3_c[4:0];
assign conv1_kernel1_3_c[0] = 16'hFCCB;
assign conv1_kernel1_3_c[1] = 16'h08BE;
assign conv1_kernel1_3_c[2] = 16'h057A;
assign conv1_kernel1_3_c[3] = 16'hFEA8;
assign conv1_kernel1_3_c[4] = 16'hFEEB;


//conv1 kernel1_4 coeff
wire signed[15:0] conv1_kernel1_4_c[4:0];
assign conv1_kernel1_4_c[0] = 16'hF899;
assign conv1_kernel1_4_c[1] = 16'h0304;
assign conv1_kernel1_4_c[2] = 16'hFA40;
assign conv1_kernel1_4_c[3] = 16'hEE94;
assign conv1_kernel1_4_c[4] = 16'h1717;


