//FC0_node0
wire signed[15:0] fc0_node0_c[29:0];
assign fc0_node0_c[0] = 16'h01F4;
assign fc0_node0_c[1] = 16'hF98C;
assign fc0_node0_c[2] = 16'hFD6A;
assign fc0_node0_c[3] = 16'h168F;
assign fc0_node0_c[4] = 16'h0568;
assign fc0_node0_c[5] = 16'hF6F1;
assign fc0_node0_c[6] = 16'h045A;
assign fc0_node0_c[7] = 16'hF0C5;
assign fc0_node0_c[8] = 16'hFB9F;
assign fc0_node0_c[9] = 16'h0000;
assign fc0_node0_c[10] = 16'h0000;
assign fc0_node0_c[11] = 16'h0000;
assign fc0_node0_c[12] = 16'h0000;
assign fc0_node0_c[13] = 16'hFDF3;
assign fc0_node0_c[14] = 16'h0000;
assign fc0_node0_c[15] = 16'h0000;
assign fc0_node0_c[16] = 16'hF383;
assign fc0_node0_c[17] = 16'hF550;
assign fc0_node0_c[18] = 16'h036E;
assign fc0_node0_c[19] = 16'h13A0;
assign fc0_node0_c[20] = 16'h0368;
assign fc0_node0_c[21] = 16'hEFD9;
assign fc0_node0_c[22] = 16'h0C52;
assign fc0_node0_c[23] = 16'h0000;
assign fc0_node0_c[24] = 16'hEE1B;
assign fc0_node0_c[25] = 16'h061C;
assign fc0_node0_c[26] = 16'h0C2D;
assign fc0_node0_c[27] = 16'h0000;
assign fc0_node0_c[28] = 16'h0766;
assign fc0_node0_c[29] = 16'hF7C7;


//FC0_node1
wire signed[15:0] fc0_node1_c[29:0];
assign fc0_node1_c[0] = 16'h025F;
assign fc0_node1_c[1] = 16'hF7C1;
assign fc0_node1_c[2] = 16'hFC74;
assign fc0_node1_c[3] = 16'h0FBB;
assign fc0_node1_c[4] = 16'h079F;
assign fc0_node1_c[5] = 16'hFD1A;
assign fc0_node1_c[6] = 16'h0288;
assign fc0_node1_c[7] = 16'hF6EE;
assign fc0_node1_c[8] = 16'h0000;
assign fc0_node1_c[9] = 16'hFD07;
assign fc0_node1_c[10] = 16'hFBED;
assign fc0_node1_c[11] = 16'h0000;
assign fc0_node1_c[12] = 16'h0000;
assign fc0_node1_c[13] = 16'hFDB8;
assign fc0_node1_c[14] = 16'h0384;
assign fc0_node1_c[15] = 16'h050C;
assign fc0_node1_c[16] = 16'hFC0C;
assign fc0_node1_c[17] = 16'h0000;
assign fc0_node1_c[18] = 16'h0000;
assign fc0_node1_c[19] = 16'h0602;
assign fc0_node1_c[20] = 16'h0000;
assign fc0_node1_c[21] = 16'hFBD3;
assign fc0_node1_c[22] = 16'h0000;
assign fc0_node1_c[23] = 16'hFC7D;
assign fc0_node1_c[24] = 16'hF094;
assign fc0_node1_c[25] = 16'h0000;
assign fc0_node1_c[26] = 16'h0811;
assign fc0_node1_c[27] = 16'h0493;
assign fc0_node1_c[28] = 16'h048E;
assign fc0_node1_c[29] = 16'h02A3;


//FC0_node2
wire signed[15:0] fc0_node2_c[29:0];
assign fc0_node2_c[0] = 16'h02E6;
assign fc0_node2_c[1] = 16'h036A;
assign fc0_node2_c[2] = 16'h0000;
assign fc0_node2_c[3] = 16'h0C64;
assign fc0_node2_c[4] = 16'h0253;
assign fc0_node2_c[5] = 16'hFB1C;
assign fc0_node2_c[6] = 16'hF9E0;
assign fc0_node2_c[7] = 16'h0484;
assign fc0_node2_c[8] = 16'h0C6C;
assign fc0_node2_c[9] = 16'hEE6D;
assign fc0_node2_c[10] = 16'h033D;
assign fc0_node2_c[11] = 16'hFDE0;
assign fc0_node2_c[12] = 16'h0000;
assign fc0_node2_c[13] = 16'hFC5A;
assign fc0_node2_c[14] = 16'h0000;
assign fc0_node2_c[15] = 16'hFDB4;
assign fc0_node2_c[16] = 16'hFA47;
assign fc0_node2_c[17] = 16'h0000;
assign fc0_node2_c[18] = 16'hF539;
assign fc0_node2_c[19] = 16'h05F3;
assign fc0_node2_c[20] = 16'h0000;
assign fc0_node2_c[21] = 16'h1362;
assign fc0_node2_c[22] = 16'hF734;
assign fc0_node2_c[23] = 16'hEE29;
assign fc0_node2_c[24] = 16'hE914;
assign fc0_node2_c[25] = 16'h0C4A;
assign fc0_node2_c[26] = 16'h0C7E;
assign fc0_node2_c[27] = 16'h0CDD;
assign fc0_node2_c[28] = 16'h16F7;
assign fc0_node2_c[29] = 16'h0000;


//FC0_node3
wire signed[15:0] fc0_node3_c[29:0];
assign fc0_node3_c[0] = 16'h04A2;
assign fc0_node3_c[1] = 16'h0000;
assign fc0_node3_c[2] = 16'h0000;
assign fc0_node3_c[3] = 16'hFDD7;
assign fc0_node3_c[4] = 16'h01AF;
assign fc0_node3_c[5] = 16'h03AF;
assign fc0_node3_c[6] = 16'hF811;
assign fc0_node3_c[7] = 16'h0AEA;
assign fc0_node3_c[8] = 16'h028E;
assign fc0_node3_c[9] = 16'hFBCE;
assign fc0_node3_c[10] = 16'h0000;
assign fc0_node3_c[11] = 16'hFDC5;
assign fc0_node3_c[12] = 16'hFBD0;
assign fc0_node3_c[13] = 16'h0200;
assign fc0_node3_c[14] = 16'hFE00;
assign fc0_node3_c[15] = 16'h048E;
assign fc0_node3_c[16] = 16'h05C9;
assign fc0_node3_c[17] = 16'h07C7;
assign fc0_node3_c[18] = 16'h0000;
assign fc0_node3_c[19] = 16'hF123;
assign fc0_node3_c[20] = 16'hF630;
assign fc0_node3_c[21] = 16'h0DD2;
assign fc0_node3_c[22] = 16'hF896;
assign fc0_node3_c[23] = 16'hFD77;
assign fc0_node3_c[24] = 16'h0405;
assign fc0_node3_c[25] = 16'h02C8;
assign fc0_node3_c[26] = 16'hFCB0;
assign fc0_node3_c[27] = 16'h0000;
assign fc0_node3_c[28] = 16'hFAAF;
assign fc0_node3_c[29] = 16'h032F;


//FC0_node4
wire signed[15:0] fc0_node4_c[29:0];
assign fc0_node4_c[0] = 16'hF771;
assign fc0_node4_c[1] = 16'h0000;
assign fc0_node4_c[2] = 16'h04C8;
assign fc0_node4_c[3] = 16'hF0ED;
assign fc0_node4_c[4] = 16'hF978;
assign fc0_node4_c[5] = 16'h068E;
assign fc0_node4_c[6] = 16'h1528;
assign fc0_node4_c[7] = 16'h0258;
assign fc0_node4_c[8] = 16'h0000;
assign fc0_node4_c[9] = 16'hF910;
assign fc0_node4_c[10] = 16'h06BB;
assign fc0_node4_c[11] = 16'h0000;
assign fc0_node4_c[12] = 16'h05BB;
assign fc0_node4_c[13] = 16'h0000;
assign fc0_node4_c[14] = 16'hFBFA;
assign fc0_node4_c[15] = 16'hF334;
assign fc0_node4_c[16] = 16'hFC79;
assign fc0_node4_c[17] = 16'h09B9;
assign fc0_node4_c[18] = 16'h0416;
assign fc0_node4_c[19] = 16'h196A;
assign fc0_node4_c[20] = 16'h1153;
assign fc0_node4_c[21] = 16'hF210;
assign fc0_node4_c[22] = 16'hFACD;
assign fc0_node4_c[23] = 16'hF6DE;
assign fc0_node4_c[24] = 16'hF788;
assign fc0_node4_c[25] = 16'h065C;
assign fc0_node4_c[26] = 16'h05F9;
assign fc0_node4_c[27] = 16'hF8A4;
assign fc0_node4_c[28] = 16'h091D;
assign fc0_node4_c[29] = 16'hFDCE;


//FC0_node5
wire signed[15:0] fc0_node5_c[29:0];
assign fc0_node5_c[0] = 16'h0451;
assign fc0_node5_c[1] = 16'hFBC4;
assign fc0_node5_c[2] = 16'hFCD0;
assign fc0_node5_c[3] = 16'hFA3D;
assign fc0_node5_c[4] = 16'h020D;
assign fc0_node5_c[5] = 16'h0771;
assign fc0_node5_c[6] = 16'h052E;
assign fc0_node5_c[7] = 16'h0681;
assign fc0_node5_c[8] = 16'h0000;
assign fc0_node5_c[9] = 16'h0000;
assign fc0_node5_c[10] = 16'hFA4F;
assign fc0_node5_c[11] = 16'h0000;
assign fc0_node5_c[12] = 16'hFE24;
assign fc0_node5_c[13] = 16'h0000;
assign fc0_node5_c[14] = 16'h0000;
assign fc0_node5_c[15] = 16'h056E;
assign fc0_node5_c[16] = 16'h0AB9;
assign fc0_node5_c[17] = 16'h0B9C;
assign fc0_node5_c[18] = 16'h0000;
assign fc0_node5_c[19] = 16'hF623;
assign fc0_node5_c[20] = 16'hF778;
assign fc0_node5_c[21] = 16'h074A;
assign fc0_node5_c[22] = 16'hF6C2;
assign fc0_node5_c[23] = 16'hF6F6;
assign fc0_node5_c[24] = 16'h02C5;
assign fc0_node5_c[25] = 16'hFA35;
assign fc0_node5_c[26] = 16'hFE04;
assign fc0_node5_c[27] = 16'h0799;
assign fc0_node5_c[28] = 16'hF7CE;
assign fc0_node5_c[29] = 16'h0460;


//FC0_node6
wire signed[15:0] fc0_node6_c[29:0];
assign fc0_node6_c[0] = 16'hFA59;
assign fc0_node6_c[1] = 16'h0523;
assign fc0_node6_c[2] = 16'h0443;
assign fc0_node6_c[3] = 16'hF079;
assign fc0_node6_c[4] = 16'hF3A7;
assign fc0_node6_c[5] = 16'hFD6A;
assign fc0_node6_c[6] = 16'h057C;
assign fc0_node6_c[7] = 16'h0811;
assign fc0_node6_c[8] = 16'h0A89;
assign fc0_node6_c[9] = 16'hF98C;
assign fc0_node6_c[10] = 16'h06A6;
assign fc0_node6_c[11] = 16'hFC86;
assign fc0_node6_c[12] = 16'h03D7;
assign fc0_node6_c[13] = 16'h03E6;
assign fc0_node6_c[14] = 16'h0000;
assign fc0_node6_c[15] = 16'hF65C;
assign fc0_node6_c[16] = 16'hFDF4;
assign fc0_node6_c[17] = 16'h0000;
assign fc0_node6_c[18] = 16'hFB38;
assign fc0_node6_c[19] = 16'h0978;
assign fc0_node6_c[20] = 16'h09A7;
assign fc0_node6_c[21] = 16'h052E;
assign fc0_node6_c[22] = 16'hF8FD;
assign fc0_node6_c[23] = 16'hEEAD;
assign fc0_node6_c[24] = 16'hFB5D;
assign fc0_node6_c[25] = 16'h07A0;
assign fc0_node6_c[26] = 16'h0497;
assign fc0_node6_c[27] = 16'h0000;
assign fc0_node6_c[28] = 16'h15BC;
assign fc0_node6_c[29] = 16'hFCB3;


//FC0_node7
wire signed[15:0] fc0_node7_c[29:0];
assign fc0_node7_c[0] = 16'h0000;
assign fc0_node7_c[1] = 16'h036E;
assign fc0_node7_c[2] = 16'h0000;
assign fc0_node7_c[3] = 16'hF6AE;
assign fc0_node7_c[4] = 16'hFA9D;
assign fc0_node7_c[5] = 16'hFD4D;
assign fc0_node7_c[6] = 16'h0000;
assign fc0_node7_c[7] = 16'h03BB;
assign fc0_node7_c[8] = 16'h0326;
assign fc0_node7_c[9] = 16'h0000;
assign fc0_node7_c[10] = 16'h0000;
assign fc0_node7_c[11] = 16'h0000;
assign fc0_node7_c[12] = 16'hFE2E;
assign fc0_node7_c[13] = 16'h02F8;
assign fc0_node7_c[14] = 16'hFE1B;
assign fc0_node7_c[15] = 16'hFB34;
assign fc0_node7_c[16] = 16'h0000;
assign fc0_node7_c[17] = 16'hFB86;
assign fc0_node7_c[18] = 16'hFBEB;
assign fc0_node7_c[19] = 16'hFE22;
assign fc0_node7_c[20] = 16'h0000;
assign fc0_node7_c[21] = 16'h03F5;
assign fc0_node7_c[22] = 16'h0000;
assign fc0_node7_c[23] = 16'h0000;
assign fc0_node7_c[24] = 16'h047E;
assign fc0_node7_c[25] = 16'h0000;
assign fc0_node7_c[26] = 16'h0000;
assign fc0_node7_c[27] = 16'h0000;
assign fc0_node7_c[28] = 16'h0363;
assign fc0_node7_c[29] = 16'h0000;


//FC0_node8
wire signed[15:0] fc0_node8_c[29:0];
assign fc0_node8_c[0] = 16'hFD99;
assign fc0_node8_c[1] = 16'h079C;
assign fc0_node8_c[2] = 16'h0251;
assign fc0_node8_c[3] = 16'hF22F;
assign fc0_node8_c[4] = 16'hF551;
assign fc0_node8_c[5] = 16'hFBCB;
assign fc0_node8_c[6] = 16'hFB8B;
assign fc0_node8_c[7] = 16'h0386;
assign fc0_node8_c[8] = 16'h04AC;
assign fc0_node8_c[9] = 16'h0469;
assign fc0_node8_c[10] = 16'h07C5;
assign fc0_node8_c[11] = 16'h0000;
assign fc0_node8_c[12] = 16'h0000;
assign fc0_node8_c[13] = 16'h032A;
assign fc0_node8_c[14] = 16'hFC03;
assign fc0_node8_c[15] = 16'hF524;
assign fc0_node8_c[16] = 16'hFC39;
assign fc0_node8_c[17] = 16'hFA0C;
assign fc0_node8_c[18] = 16'hFB86;
assign fc0_node8_c[19] = 16'hFB21;
assign fc0_node8_c[20] = 16'h0662;
assign fc0_node8_c[21] = 16'h0805;
assign fc0_node8_c[22] = 16'h03E7;
assign fc0_node8_c[23] = 16'h0401;
assign fc0_node8_c[24] = 16'h07A6;
assign fc0_node8_c[25] = 16'h0000;
assign fc0_node8_c[26] = 16'hFA41;
assign fc0_node8_c[27] = 16'hFA87;
assign fc0_node8_c[28] = 16'h0766;
assign fc0_node8_c[29] = 16'hF8FF;


//FC1_node0
wire signed[15:0] fc1_node0_c[8:0];
assign fc1_node0_c[0] = 16'h15A5;
assign fc1_node0_c[1] = 16'h0748;
assign fc1_node0_c[2] = 16'h0000;
assign fc1_node0_c[3] = 16'hF26A;
assign fc1_node0_c[4] = 16'h0E8E;
assign fc1_node0_c[5] = 16'hF1D4;
assign fc1_node0_c[6] = 16'h02A9;
assign fc1_node0_c[7] = 16'hFC1D;
assign fc1_node0_c[8] = 16'h0000;


//FC1_node1
wire signed[15:0] fc1_node1_c[8:0];
assign fc1_node1_c[0] = 16'h0666;
assign fc1_node1_c[1] = 16'h03B1;
assign fc1_node1_c[2] = 16'hED4F;
assign fc1_node1_c[3] = 16'hFDEC;
assign fc1_node1_c[4] = 16'hF0CD;
assign fc1_node1_c[5] = 16'h0000;
assign fc1_node1_c[6] = 16'hEB4F;
assign fc1_node1_c[7] = 16'hFB17;
assign fc1_node1_c[8] = 16'hFC98;


//FC1_node2
wire signed[15:0] fc1_node2_c[8:0];
assign fc1_node2_c[0] = 16'hFA7C;
assign fc1_node2_c[1] = 16'h0000;
assign fc1_node2_c[2] = 16'h1274;
assign fc1_node2_c[3] = 16'h05D9;
assign fc1_node2_c[4] = 16'hF224;
assign fc1_node2_c[5] = 16'h0000;
assign fc1_node2_c[6] = 16'h0B68;
assign fc1_node2_c[7] = 16'h042A;
assign fc1_node2_c[8] = 16'h0B44;


//FC1_node3
wire signed[15:0] fc1_node3_c[8:0];
assign fc1_node3_c[0] = 16'hED24;
assign fc1_node3_c[1] = 16'hF1B7;
assign fc1_node3_c[2] = 16'hEF3B;
assign fc1_node3_c[3] = 16'h04D3;
assign fc1_node3_c[4] = 16'h08A2;
assign fc1_node3_c[5] = 16'h0498;
assign fc1_node3_c[6] = 16'h0744;
assign fc1_node3_c[7] = 16'h0404;
assign fc1_node3_c[8] = 16'h0C01;


//FC1_node4
wire signed[15:0] fc1_node4_c[8:0];
assign fc1_node4_c[0] = 16'h0000;
assign fc1_node4_c[1] = 16'h0B9D;
assign fc1_node4_c[2] = 16'h171F;
assign fc1_node4_c[3] = 16'h0740;
assign fc1_node4_c[4] = 16'h08A1;
assign fc1_node4_c[5] = 16'h0C88;
assign fc1_node4_c[6] = 16'h062E;
assign fc1_node4_c[7] = 16'hF931;
assign fc1_node4_c[8] = 16'hF354;


