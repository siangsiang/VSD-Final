wire [31:0] FIR_C [99:0];
assign FIR_C[0] = 31'h0000B203;    // 0.00016976520419120789
assign FIR_C[1] = 31'h00003181;    // 0.00004721060395240784
assign FIR_C[2] = 31'hFFFF864B;    // -0.00011606886982917786
assign FIR_C[3] = 31'hFFFED465;    // -0.00028572604060173035
assign FIR_C[4] = 31'hFFFEE129;    // -0.00027355179190635681
assign FIR_C[5] = 31'h000008F9;    // 0.00000855699181556702
assign FIR_C[6] = 31'h0001A798;    // 0.00040397047996520996
assign FIR_C[7] = 31'h00024FF6;    // 0.00056453794240951538
assign FIR_C[8] = 31'h0000F1CA;    // 0.00023058801889419556
assign FIR_C[9] = 31'hFFFE1436;    // -0.00046900659799575806
assign FIR_C[10] = 31'hFFFBEE58;    // -0.00099340081214904785
assign FIR_C[11] = 31'hFFFCD644;    // -0.00077222287654876709
assign FIR_C[12] = 31'h0001036E;    // 0.00024741142988204956
assign FIR_C[13] = 31'h00059FCA;    // 0.00137308984994888306
assign FIR_C[14] = 31'h00067ED1;    // 0.00158578529953956604
assign FIR_C[15] = 31'h0001A7AB;    // 0.00040404126048088074
assign FIR_C[16] = 31'hFFF9DBAF;    // -0.00149947777390480042
assign FIR_C[17] = 31'hFFF566C7;    // -0.00258753076195716858
assign FIR_C[18] = 31'hFFF949BF;    // -0.00163865461945533752
assign FIR_C[19] = 31'h000442E3;    // 0.00104035064578056335
assign FIR_C[20] = 31'h000E4861;    // 0.00348699465394020081
assign FIR_C[21] = 31'h000E18D4;    // 0.00344164669513702393
assign FIR_C[22] = 31'h00015094;    // 0.00032098591327667236
assign FIR_C[23] = 31'hFFF04341;    // -0.00384211167693138123
assign FIR_C[24] = 31'hFFE91589;    // -0.00559469684958457947
assign FIR_C[25] = 31'hFFF4752F;    // -0.00281793251633644104
assign FIR_C[26] = 31'h000C9948;    // 0.00307586789131164551
assign FIR_C[27] = 31'h001F1C74;    // 0.00759549438953399658
assign FIR_C[28] = 31'h001A729E;    // 0.00645696371793746948
assign FIR_C[29] = 31'hFFFD943B;    // -0.00059105828404426575
assign FIR_C[30] = 31'hFFDC8104;    // -0.00866602361202239990
assign FIR_C[31] = 31'hFFD342CF;    // -0.01092261448502540588
assign FIR_C[32] = 31'hFFEF2149;    // -0.00411864742636680603
assign FIR_C[33] = 31'h001FDF2C;    // 0.00778119266033172607
assign FIR_C[34] = 31'h003F8169;    // 0.01550427451729774475
assign FIR_C[35] = 31'h002E9588;    // 0.01137307286262512207
assign FIR_C[36] = 31'hFFF0DF30;    // -0.00369340181350708008
assign FIR_C[37] = 31'hFFB1ED1B;    // -0.01906098797917366028
assign FIR_C[38] = 31'hFFA89835;    // -0.02133921906352043152
assign FIR_C[39] = 31'hFFEA81BB;    // -0.00524737313389778137
assign FIR_C[40] = 31'h00517CAA;    // 0.01989427953958511353
assign FIR_C[41] = 31'h008CEDEC;    // 0.03440658748149871826
assign FIR_C[42] = 31'h005AB35B;    // 0.02214370295405387878
assign FIR_C[43] = 31'hFFC2B5A1;    // -0.01496350392699241638
assign FIR_C[44] = 31'hFF272F92;    // -0.05293314903974533081
assign FIR_C[45] = 31'hFF147F7A;    // -0.05749561637639999390
assign FIR_C[46] = 31'hFFE7CF85;    // -0.00590560957789421082
assign FIR_C[47] = 31'h01853667;    // 0.09502258524298667908
assign FIR_C[48] = 31'h035259BC;    // 0.20760510861873626709
assign FIR_C[49] = 31'h04812148;    // 0.28152588009834289551
assign FIR_C[50] = 31'h04812148;    // 0.28152588009834289551
assign FIR_C[51] = 31'h035259BC;    // 0.20760510861873626709
assign FIR_C[52] = 31'h01853667;    // 0.09502258524298667908
assign FIR_C[53] = 31'hFFE7CF85;    // -0.00590560957789421082
assign FIR_C[54] = 31'hFF147F7A;    // -0.05749561637639999390
assign FIR_C[55] = 31'hFF272F92;    // -0.05293314903974533081
assign FIR_C[56] = 31'hFFC2B5A1;    // -0.01496350392699241638
assign FIR_C[57] = 31'h005AB35B;    // 0.02214370295405387878
assign FIR_C[58] = 31'h008CEDEC;    // 0.03440658748149871826
assign FIR_C[59] = 31'h00517CAA;    // 0.01989427953958511353
assign FIR_C[60] = 31'hFFEA81BB;    // -0.00524737313389778137
assign FIR_C[61] = 31'hFFA89835;    // -0.02133921906352043152
assign FIR_C[62] = 31'hFFB1ED1B;    // -0.01906098797917366028
assign FIR_C[63] = 31'hFFF0DF30;    // -0.00369340181350708008
assign FIR_C[64] = 31'h002E9588;    // 0.01137307286262512207
assign FIR_C[65] = 31'h003F8169;    // 0.01550427451729774475
assign FIR_C[66] = 31'h001FDF2C;    // 0.00778119266033172607
assign FIR_C[67] = 31'hFFEF2149;    // -0.00411864742636680603
assign FIR_C[68] = 31'hFFD342CF;    // -0.01092261448502540588
assign FIR_C[69] = 31'hFFDC8104;    // -0.00866602361202239990
assign FIR_C[70] = 31'hFFFD943B;    // -0.00059105828404426575
assign FIR_C[71] = 31'h001A729E;    // 0.00645696371793746948
assign FIR_C[72] = 31'h001F1C74;    // 0.00759549438953399658
assign FIR_C[73] = 31'h000C9948;    // 0.00307586789131164551
assign FIR_C[74] = 31'hFFF4752F;    // -0.00281793251633644104
assign FIR_C[75] = 31'hFFE91589;    // -0.00559469684958457947
assign FIR_C[76] = 31'hFFF04341;    // -0.00384211167693138123
assign FIR_C[77] = 31'h00015094;    // 0.00032098591327667236
assign FIR_C[78] = 31'h000E18D4;    // 0.00344164669513702393
assign FIR_C[79] = 31'h000E4861;    // 0.00348699465394020081
assign FIR_C[80] = 31'h000442E3;    // 0.00104035064578056335
assign FIR_C[81] = 31'hFFF949BF;    // -0.00163865461945533752
assign FIR_C[82] = 31'hFFF566C7;    // -0.00258753076195716858
assign FIR_C[83] = 31'hFFF9DBAF;    // -0.00149947777390480042
assign FIR_C[84] = 31'h0001A7AB;    // 0.00040404126048088074
assign FIR_C[85] = 31'h00067ED1;    // 0.00158578529953956604
assign FIR_C[86] = 31'h00059FCA;    // 0.00137308984994888306
assign FIR_C[87] = 31'h0001036E;    // 0.00024741142988204956
assign FIR_C[88] = 31'hFFFCD644;    // -0.00077222287654876709
assign FIR_C[89] = 31'hFFFBEE58;    // -0.00099340081214904785
assign FIR_C[90] = 31'hFFFE1436;    // -0.00046900659799575806
assign FIR_C[91] = 31'h0000F1CA;    // 0.00023058801889419556
assign FIR_C[92] = 31'h00024FF6;    // 0.00056453794240951538
assign FIR_C[93] = 31'h0001A798;    // 0.00040397047996520996
assign FIR_C[94] = 31'h000008F9;    // 0.00000855699181556702
assign FIR_C[95] = 31'hFFFEE129;    // -0.00027355179190635681
assign FIR_C[96] = 31'hFFFED465;    // -0.00028572604060173035
assign FIR_C[97] = 31'hFFFF864B;    // -0.00011606886982917786
assign FIR_C[98] = 31'h00003181;    // 0.00004721060395240784
assign FIR_C[99] = 31'h0000B203;    // 0.00016976520419120789
