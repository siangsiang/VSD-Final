reg [15:0] FIR_C0 = 16'h0000;    // 0.00000000000000000000
reg [15:0] FIR_C1 = 16'h0000;    // 0.00000000000000000000
reg [15:0] FIR_C2 = 16'h0000;    // 0.00000000000000000000
reg [15:0] FIR_C3 = 16'hFFFF;    // -0.00024414062500000000
reg [15:0] FIR_C4 = 16'hFFFF;    // -0.00024414062500000000
reg [15:0] FIR_C5 = 16'h0000;    // 0.00000000000000000000
reg [15:0] FIR_C6 = 16'h0001;    // 0.00024414062500000000
reg [15:0] FIR_C7 = 16'h0002;    // 0.00048828125000000000
reg [15:0] FIR_C8 = 16'h0000;    // 0.00000000000000000000
reg [15:0] FIR_C9 = 16'hFFFF;    // -0.00024414062500000000
reg [15:0] FIR_C10 = 16'hFFFC;    // -0.00097656250000000000
reg [15:0] FIR_C11 = 16'hFFFD;    // -0.00073242187500000000
reg [15:0] FIR_C12 = 16'h0001;    // 0.00024414062500000000
reg [15:0] FIR_C13 = 16'h0005;    // 0.00122070312500000000
reg [15:0] FIR_C14 = 16'h0006;    // 0.00146484375000000000
reg [15:0] FIR_C15 = 16'h0001;    // 0.00024414062500000000
reg [15:0] FIR_C16 = 16'hFFFA;    // -0.00146484375000000000
reg [15:0] FIR_C17 = 16'hFFF6;    // -0.00244140625000000000
reg [15:0] FIR_C18 = 16'hFFFA;    // -0.00146484375000000000
reg [15:0] FIR_C19 = 16'h0004;    // 0.00097656250000000000
reg [15:0] FIR_C20 = 16'h000E;    // 0.00341796875000000000
reg [15:0] FIR_C21 = 16'h000E;    // 0.00341796875000000000
reg [15:0] FIR_C22 = 16'h0001;    // 0.00024414062500000000
reg [15:0] FIR_C23 = 16'hFFF1;    // -0.00366210937500000000
reg [15:0] FIR_C24 = 16'hFFEA;    // -0.00537109375000000000
reg [15:0] FIR_C25 = 16'hFFF5;    // -0.00268554687500000000
reg [15:0] FIR_C26 = 16'h000C;    // 0.00292968750000000000
reg [15:0] FIR_C27 = 16'h001F;    // 0.00756835937500000000
reg [15:0] FIR_C28 = 16'h001A;    // 0.00634765625000000000
reg [15:0] FIR_C29 = 16'hFFFE;    // -0.00048828125000000000
reg [15:0] FIR_C30 = 16'hFFDD;    // -0.00854492187500000000
reg [15:0] FIR_C31 = 16'hFFD4;    // -0.01074218750000000000
reg [15:0] FIR_C32 = 16'hFFF0;    // -0.00390625000000000000
reg [15:0] FIR_C33 = 16'h001F;    // 0.00756835937500000000
reg [15:0] FIR_C34 = 16'h003F;    // 0.01538085937500000000
reg [15:0] FIR_C35 = 16'h002E;    // 0.01123046875000000000
reg [15:0] FIR_C36 = 16'hFFF1;    // -0.00366210937500000000
reg [15:0] FIR_C37 = 16'hFFB2;    // -0.01904296875000000000
reg [15:0] FIR_C38 = 16'hFFA9;    // -0.02124023437500000000
reg [15:0] FIR_C39 = 16'hFFEB;    // -0.00512695312500000000
reg [15:0] FIR_C40 = 16'h0051;    // 0.01977539062500000000
reg [15:0] FIR_C41 = 16'h008C;    // 0.03417968750000000000
reg [15:0] FIR_C42 = 16'h005A;    // 0.02197265625000000000
reg [15:0] FIR_C43 = 16'hFFC3;    // -0.01489257812500000000
reg [15:0] FIR_C44 = 16'hFF28;    // -0.05273437500000000000
reg [15:0] FIR_C45 = 16'hFF15;    // -0.05737304687500000000
reg [15:0] FIR_C46 = 16'hFFE8;    // -0.00585937500000000000
reg [15:0] FIR_C47 = 16'h0185;    // 0.09497070312500000000
reg [15:0] FIR_C48 = 16'h0352;    // 0.20751953125000000000
reg [15:0] FIR_C49 = 16'h0481;    // 0.28149414062500000000
reg [15:0] FIR_C50 = 16'h0481;    // 0.28149414062500000000
reg [15:0] FIR_C51 = 16'h0352;    // 0.20751953125000000000
reg [15:0] FIR_C52 = 16'h0185;    // 0.09497070312500000000
reg [15:0] FIR_C53 = 16'hFFE8;    // -0.00585937500000000000
reg [15:0] FIR_C54 = 16'hFF15;    // -0.05737304687500000000
reg [15:0] FIR_C55 = 16'hFF28;    // -0.05273437500000000000
reg [15:0] FIR_C56 = 16'hFFC3;    // -0.01489257812500000000
reg [15:0] FIR_C57 = 16'h005A;    // 0.02197265625000000000
reg [15:0] FIR_C58 = 16'h008C;    // 0.03417968750000000000
reg [15:0] FIR_C59 = 16'h0051;    // 0.01977539062500000000
reg [15:0] FIR_C60 = 16'hFFEB;    // -0.00512695312500000000
reg [15:0] FIR_C61 = 16'hFFA9;    // -0.02124023437500000000
reg [15:0] FIR_C62 = 16'hFFB2;    // -0.01904296875000000000
reg [15:0] FIR_C63 = 16'hFFF1;    // -0.00366210937500000000
reg [15:0] FIR_C64 = 16'h002E;    // 0.01123046875000000000
reg [15:0] FIR_C65 = 16'h003F;    // 0.01538085937500000000
reg [15:0] FIR_C66 = 16'h001F;    // 0.00756835937500000000
reg [15:0] FIR_C67 = 16'hFFF0;    // -0.00390625000000000000
reg [15:0] FIR_C68 = 16'hFFD4;    // -0.01074218750000000000
reg [15:0] FIR_C69 = 16'hFFDD;    // -0.00854492187500000000
reg [15:0] FIR_C70 = 16'hFFFE;    // -0.00048828125000000000
reg [15:0] FIR_C71 = 16'h001A;    // 0.00634765625000000000
reg [15:0] FIR_C72 = 16'h001F;    // 0.00756835937500000000
reg [15:0] FIR_C73 = 16'h000C;    // 0.00292968750000000000
reg [15:0] FIR_C74 = 16'hFFF5;    // -0.00268554687500000000
reg [15:0] FIR_C75 = 16'hFFEA;    // -0.00537109375000000000
reg [15:0] FIR_C76 = 16'hFFF1;    // -0.00366210937500000000
reg [15:0] FIR_C77 = 16'h0001;    // 0.00024414062500000000
reg [15:0] FIR_C78 = 16'h000E;    // 0.00341796875000000000
reg [15:0] FIR_C79 = 16'h000E;    // 0.00341796875000000000
reg [15:0] FIR_C80 = 16'h0004;    // 0.00097656250000000000
reg [15:0] FIR_C81 = 16'hFFFA;    // -0.00146484375000000000
reg [15:0] FIR_C82 = 16'hFFF6;    // -0.00244140625000000000
reg [15:0] FIR_C83 = 16'hFFFA;    // -0.00146484375000000000
reg [15:0] FIR_C84 = 16'h0001;    // 0.00024414062500000000
reg [15:0] FIR_C85 = 16'h0006;    // 0.00146484375000000000
reg [15:0] FIR_C86 = 16'h0005;    // 0.00122070312500000000
reg [15:0] FIR_C87 = 16'h0001;    // 0.00024414062500000000
reg [15:0] FIR_C88 = 16'hFFFD;    // -0.00073242187500000000
reg [15:0] FIR_C89 = 16'hFFFC;    // -0.00097656250000000000
reg [15:0] FIR_C90 = 16'hFFFF;    // -0.00024414062500000000
reg [15:0] FIR_C91 = 16'h0000;    // 0.00000000000000000000
reg [15:0] FIR_C92 = 16'h0002;    // 0.00048828125000000000
reg [15:0] FIR_C93 = 16'h0001;    // 0.00024414062500000000
reg [15:0] FIR_C94 = 16'h0000;    // 0.00000000000000000000
reg [15:0] FIR_C95 = 16'hFFFF;    // -0.00024414062500000000
reg [15:0] FIR_C96 = 16'hFFFF;    // -0.00024414062500000000
reg [15:0] FIR_C97 = 16'h0000;    // 0.00000000000000000000
reg [15:0] FIR_C98 = 16'h0000;    // 0.00000000000000000000
reg [15:0] FIR_C99 = 16'h0000;    // 0.00000000000000000000
