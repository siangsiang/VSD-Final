//FC0_node0
wire signed[15:0] fc0_node0_c[29:0];
assign fc0_node0_c[0] = 16'h07DA;
assign fc0_node0_c[1] = 16'hF660;
assign fc0_node0_c[2] = 16'hFCA0;
assign fc0_node0_c[3] = 16'h1910;
assign fc0_node0_c[4] = 16'h0059;
assign fc0_node0_c[5] = 16'hF669;
assign fc0_node0_c[6] = 16'h0205;
assign fc0_node0_c[7] = 16'hF642;
assign fc0_node0_c[8] = 16'hF972;
assign fc0_node0_c[9] = 16'h01A6;
assign fc0_node0_c[10] = 16'h03F8;
assign fc0_node0_c[11] = 16'hFEAF;
assign fc0_node0_c[12] = 16'hFEA6;
assign fc0_node0_c[13] = 16'h0072;
assign fc0_node0_c[14] = 16'hFF89;
assign fc0_node0_c[15] = 16'h0207;
assign fc0_node0_c[16] = 16'hF41B;
assign fc0_node0_c[17] = 16'hF896;
assign fc0_node0_c[18] = 16'hFD60;
assign fc0_node0_c[19] = 16'h105B;
assign fc0_node0_c[20] = 16'h0438;
assign fc0_node0_c[21] = 16'hEED3;
assign fc0_node0_c[22] = 16'h0A35;
assign fc0_node0_c[23] = 16'hFD2A;
assign fc0_node0_c[24] = 16'hEFB7;
assign fc0_node0_c[25] = 16'h0627;
assign fc0_node0_c[26] = 16'h0BDB;
assign fc0_node0_c[27] = 16'h037D;
assign fc0_node0_c[28] = 16'h09EE;
assign fc0_node0_c[29] = 16'hF871;


//FC0_node1
wire signed[15:0] fc0_node1_c[29:0];
assign fc0_node1_c[0] = 16'h04F4;
assign fc0_node1_c[1] = 16'hF772;
assign fc0_node1_c[2] = 16'hFCBA;
assign fc0_node1_c[3] = 16'h109D;
assign fc0_node1_c[4] = 16'h0301;
assign fc0_node1_c[5] = 16'hFC62;
assign fc0_node1_c[6] = 16'h019D;
assign fc0_node1_c[7] = 16'hFB99;
assign fc0_node1_c[8] = 16'hFF07;
assign fc0_node1_c[9] = 16'hFF08;
assign fc0_node1_c[10] = 16'hFD2C;
assign fc0_node1_c[11] = 16'h001D;
assign fc0_node1_c[12] = 16'h01FE;
assign fc0_node1_c[13] = 16'hFE8E;
assign fc0_node1_c[14] = 16'h01E6;
assign fc0_node1_c[15] = 16'h0548;
assign fc0_node1_c[16] = 16'hFB9C;
assign fc0_node1_c[17] = 16'hFE3D;
assign fc0_node1_c[18] = 16'hFF5B;
assign fc0_node1_c[19] = 16'h076E;
assign fc0_node1_c[20] = 16'hFF37;
assign fc0_node1_c[21] = 16'hFA7D;
assign fc0_node1_c[22] = 16'h0028;
assign fc0_node1_c[23] = 16'hFE14;
assign fc0_node1_c[24] = 16'hF3CF;
assign fc0_node1_c[25] = 16'h009E;
assign fc0_node1_c[26] = 16'h0743;
assign fc0_node1_c[27] = 16'h03A5;
assign fc0_node1_c[28] = 16'h04A3;
assign fc0_node1_c[29] = 16'h020E;


//FC0_node2
wire signed[15:0] fc0_node2_c[29:0];
assign fc0_node2_c[0] = 16'h0675;
assign fc0_node2_c[1] = 16'h0299;
assign fc0_node2_c[2] = 16'h024E;
assign fc0_node2_c[3] = 16'h0D31;
assign fc0_node2_c[4] = 16'hFB4F;
assign fc0_node2_c[5] = 16'hF92F;
assign fc0_node2_c[6] = 16'hFD68;
assign fc0_node2_c[7] = 16'h05C2;
assign fc0_node2_c[8] = 16'h06F4;
assign fc0_node2_c[9] = 16'hF233;
assign fc0_node2_c[10] = 16'h0172;
assign fc0_node2_c[11] = 16'h0118;
assign fc0_node2_c[12] = 16'h03EA;
assign fc0_node2_c[13] = 16'hFD8C;
assign fc0_node2_c[14] = 16'hFF4A;
assign fc0_node2_c[15] = 16'h020E;
assign fc0_node2_c[16] = 16'hF9C3;
assign fc0_node2_c[17] = 16'h0042;
assign fc0_node2_c[18] = 16'hF514;
assign fc0_node2_c[19] = 16'h079E;
assign fc0_node2_c[20] = 16'h0244;
assign fc0_node2_c[21] = 16'h14B5;
assign fc0_node2_c[22] = 16'hF4D6;
assign fc0_node2_c[23] = 16'hF24D;
assign fc0_node2_c[24] = 16'hEDD3;
assign fc0_node2_c[25] = 16'h0BE2;
assign fc0_node2_c[26] = 16'h0E91;
assign fc0_node2_c[27] = 16'h05B9;
assign fc0_node2_c[28] = 16'h1362;
assign fc0_node2_c[29] = 16'hFC2D;


//FC0_node3
wire signed[15:0] fc0_node3_c[29:0];
assign fc0_node3_c[0] = 16'h01B8;
assign fc0_node3_c[1] = 16'h0324;
assign fc0_node3_c[2] = 16'h02F6;
assign fc0_node3_c[3] = 16'hFCD6;
assign fc0_node3_c[4] = 16'h01CF;
assign fc0_node3_c[5] = 16'h0337;
assign fc0_node3_c[6] = 16'hFA27;
assign fc0_node3_c[7] = 16'h09B7;
assign fc0_node3_c[8] = 16'h024A;
assign fc0_node3_c[9] = 16'hFA83;
assign fc0_node3_c[10] = 16'hFD27;
assign fc0_node3_c[11] = 16'h0021;
assign fc0_node3_c[12] = 16'hFE1B;
assign fc0_node3_c[13] = 16'h0099;
assign fc0_node3_c[14] = 16'hFEBD;
assign fc0_node3_c[15] = 16'h0431;
assign fc0_node3_c[16] = 16'h05FE;
assign fc0_node3_c[17] = 16'h0679;
assign fc0_node3_c[18] = 16'h0328;
assign fc0_node3_c[19] = 16'hF431;
assign fc0_node3_c[20] = 16'hF4F2;
assign fc0_node3_c[21] = 16'h0F65;
assign fc0_node3_c[22] = 16'hF8F8;
assign fc0_node3_c[23] = 16'h01CC;
assign fc0_node3_c[24] = 16'h046F;
assign fc0_node3_c[25] = 16'h0238;
assign fc0_node3_c[26] = 16'hFD7B;
assign fc0_node3_c[27] = 16'hFD32;
assign fc0_node3_c[28] = 16'hF9E0;
assign fc0_node3_c[29] = 16'h0210;


//FC0_node4
wire signed[15:0] fc0_node4_c[29:0];
assign fc0_node4_c[0] = 16'hFCBA;
assign fc0_node4_c[1] = 16'hFE76;
assign fc0_node4_c[2] = 16'h00A9;
assign fc0_node4_c[3] = 16'hF167;
assign fc0_node4_c[4] = 16'hFAAE;
assign fc0_node4_c[5] = 16'h091C;
assign fc0_node4_c[6] = 16'h1334;
assign fc0_node4_c[7] = 16'h03C1;
assign fc0_node4_c[8] = 16'hFD1F;
assign fc0_node4_c[9] = 16'hFD13;
assign fc0_node4_c[10] = 16'h06A6;
assign fc0_node4_c[11] = 16'hFC08;
assign fc0_node4_c[12] = 16'h063C;
assign fc0_node4_c[13] = 16'h0037;
assign fc0_node4_c[14] = 16'hF8A7;
assign fc0_node4_c[15] = 16'hF17A;
assign fc0_node4_c[16] = 16'hF6A4;
assign fc0_node4_c[17] = 16'h06C7;
assign fc0_node4_c[18] = 16'h0618;
assign fc0_node4_c[19] = 16'h1AD8;
assign fc0_node4_c[20] = 16'h14DD;
assign fc0_node4_c[21] = 16'hEE1C;
assign fc0_node4_c[22] = 16'hFCC4;
assign fc0_node4_c[23] = 16'hF3F0;
assign fc0_node4_c[24] = 16'hF8FE;
assign fc0_node4_c[25] = 16'h05C7;
assign fc0_node4_c[26] = 16'h04F7;
assign fc0_node4_c[27] = 16'hFA46;
assign fc0_node4_c[28] = 16'h0792;
assign fc0_node4_c[29] = 16'hFE9B;


//FC0_node5
wire signed[15:0] fc0_node5_c[29:0];
assign fc0_node5_c[0] = 16'h021F;
assign fc0_node5_c[1] = 16'hFF3D;
assign fc0_node5_c[2] = 16'hFDE0;
assign fc0_node5_c[3] = 16'hFAF8;
assign fc0_node5_c[4] = 16'h0167;
assign fc0_node5_c[5] = 16'h0579;
assign fc0_node5_c[6] = 16'h0439;
assign fc0_node5_c[7] = 16'h06C1;
assign fc0_node5_c[8] = 16'h018F;
assign fc0_node5_c[9] = 16'hFDB6;
assign fc0_node5_c[10] = 16'hF919;
assign fc0_node5_c[11] = 16'h040D;
assign fc0_node5_c[12] = 16'h01BF;
assign fc0_node5_c[13] = 16'hFE40;
assign fc0_node5_c[14] = 16'h01A2;
assign fc0_node5_c[15] = 16'h051B;
assign fc0_node5_c[16] = 16'h0947;
assign fc0_node5_c[17] = 16'h0751;
assign fc0_node5_c[18] = 16'h018A;
assign fc0_node5_c[19] = 16'hFC29;
assign fc0_node5_c[20] = 16'hF7D0;
assign fc0_node5_c[21] = 16'h09D6;
assign fc0_node5_c[22] = 16'hF6AA;
assign fc0_node5_c[23] = 16'hFA79;
assign fc0_node5_c[24] = 16'h02D2;
assign fc0_node5_c[25] = 16'hFA4A;
assign fc0_node5_c[26] = 16'hFF61;
assign fc0_node5_c[27] = 16'h0573;
assign fc0_node5_c[28] = 16'hF914;
assign fc0_node5_c[29] = 16'h0320;


//FC0_node6
wire signed[15:0] fc0_node6_c[29:0];
assign fc0_node6_c[0] = 16'hFC8B;
assign fc0_node6_c[1] = 16'h0355;
assign fc0_node6_c[2] = 16'h02DC;
assign fc0_node6_c[3] = 16'hF14C;
assign fc0_node6_c[4] = 16'hF383;
assign fc0_node6_c[5] = 16'hFC0F;
assign fc0_node6_c[6] = 16'h065A;
assign fc0_node6_c[7] = 16'h0458;
assign fc0_node6_c[8] = 16'h09F0;
assign fc0_node6_c[9] = 16'hFB9F;
assign fc0_node6_c[10] = 16'h0573;
assign fc0_node6_c[11] = 16'hFCA0;
assign fc0_node6_c[12] = 16'h03F8;
assign fc0_node6_c[13] = 16'h0592;
assign fc0_node6_c[14] = 16'hFE36;
assign fc0_node6_c[15] = 16'hF9C5;
assign fc0_node6_c[16] = 16'hFBD4;
assign fc0_node6_c[17] = 16'h004E;
assign fc0_node6_c[18] = 16'hFC6F;
assign fc0_node6_c[19] = 16'h07D9;
assign fc0_node6_c[20] = 16'h0DF7;
assign fc0_node6_c[21] = 16'h06C5;
assign fc0_node6_c[22] = 16'hF87D;
assign fc0_node6_c[23] = 16'hED88;
assign fc0_node6_c[24] = 16'hFB32;
assign fc0_node6_c[25] = 16'h0834;
assign fc0_node6_c[26] = 16'h072B;
assign fc0_node6_c[27] = 16'hFED5;
assign fc0_node6_c[28] = 16'h13B1;
assign fc0_node6_c[29] = 16'hFAF0;


//FC0_node7
wire signed[15:0] fc0_node7_c[29:0];
assign fc0_node7_c[0] = 16'hFF65;
assign fc0_node7_c[1] = 16'h0365;
assign fc0_node7_c[2] = 16'h01A5;
assign fc0_node7_c[3] = 16'hF5DC;
assign fc0_node7_c[4] = 16'hFB98;
assign fc0_node7_c[5] = 16'hFC6E;
assign fc0_node7_c[6] = 16'hFFF2;
assign fc0_node7_c[7] = 16'h0061;
assign fc0_node7_c[8] = 16'h04E6;
assign fc0_node7_c[9] = 16'hFFE7;
assign fc0_node7_c[10] = 16'h00CD;
assign fc0_node7_c[11] = 16'h014A;
assign fc0_node7_c[12] = 16'hFD30;
assign fc0_node7_c[13] = 16'h036C;
assign fc0_node7_c[14] = 16'hFF02;
assign fc0_node7_c[15] = 16'hFC99;
assign fc0_node7_c[16] = 16'h0201;
assign fc0_node7_c[17] = 16'hFC35;
assign fc0_node7_c[18] = 16'hFC1B;
assign fc0_node7_c[19] = 16'hFC75;
assign fc0_node7_c[20] = 16'h029F;
assign fc0_node7_c[21] = 16'h05BC;
assign fc0_node7_c[22] = 16'hFFAF;
assign fc0_node7_c[23] = 16'hFDC2;
assign fc0_node7_c[24] = 16'h02F6;
assign fc0_node7_c[25] = 16'hFFB1;
assign fc0_node7_c[26] = 16'h006C;
assign fc0_node7_c[27] = 16'h0038;
assign fc0_node7_c[28] = 16'h03E4;
assign fc0_node7_c[29] = 16'hFED1;


//FC0_node8
wire signed[15:0] fc0_node8_c[29:0];
assign fc0_node8_c[0] = 16'hFB6E;
assign fc0_node8_c[1] = 16'h0684;
assign fc0_node8_c[2] = 16'h0211;
assign fc0_node8_c[3] = 16'hEF07;
assign fc0_node8_c[4] = 16'hF81E;
assign fc0_node8_c[5] = 16'hFBB9;
assign fc0_node8_c[6] = 16'hFD97;
assign fc0_node8_c[7] = 16'hFD70;
assign fc0_node8_c[8] = 16'h07A0;
assign fc0_node8_c[9] = 16'h042E;
assign fc0_node8_c[10] = 16'h07ED;
assign fc0_node8_c[11] = 16'hFE2E;
assign fc0_node8_c[12] = 16'hFBFA;
assign fc0_node8_c[13] = 16'h047E;
assign fc0_node8_c[14] = 16'hFD3E;
assign fc0_node8_c[15] = 16'hF6DC;
assign fc0_node8_c[16] = 16'hFDED;
assign fc0_node8_c[17] = 16'hFCD5;
assign fc0_node8_c[18] = 16'hFC9F;
assign fc0_node8_c[19] = 16'hF5FA;
assign fc0_node8_c[20] = 16'h0881;
assign fc0_node8_c[21] = 16'h08E0;
assign fc0_node8_c[22] = 16'h03A2;
assign fc0_node8_c[23] = 16'h00C4;
assign fc0_node8_c[24] = 16'h0562;
assign fc0_node8_c[25] = 16'h0341;
assign fc0_node8_c[26] = 16'hFB98;
assign fc0_node8_c[27] = 16'hFAD5;
assign fc0_node8_c[28] = 16'h06EB;
assign fc0_node8_c[29] = 16'hF881;


//FC1_node0
wire signed[15:0] fc1_node0_c[8:0];
assign fc1_node0_c[0] = 16'h153A;
assign fc1_node0_c[1] = 16'h088B;
assign fc1_node0_c[2] = 16'hFF5F;
assign fc1_node0_c[3] = 16'hF329;
assign fc1_node0_c[4] = 16'h0DF2;
assign fc1_node0_c[5] = 16'hF44B;
assign fc1_node0_c[6] = 16'h026E;
assign fc1_node0_c[7] = 16'hFB9E;
assign fc1_node0_c[8] = 16'h00AD;


//FC1_node1
wire signed[15:0] fc1_node1_c[8:0];
assign fc1_node1_c[0] = 16'h01DA;
assign fc1_node1_c[1] = 16'h022C;
assign fc1_node1_c[2] = 16'hEF56;
assign fc1_node1_c[3] = 16'hFFC0;
assign fc1_node1_c[4] = 16'hEFD7;
assign fc1_node1_c[5] = 16'hFF42;
assign fc1_node1_c[6] = 16'hEC85;
assign fc1_node1_c[7] = 16'hFB13;
assign fc1_node1_c[8] = 16'hFD4C;


//FC1_node2
wire signed[15:0] fc1_node2_c[8:0];
assign fc1_node2_c[0] = 16'hFD0C;
assign fc1_node2_c[1] = 16'h001B;
assign fc1_node2_c[2] = 16'h11E2;
assign fc1_node2_c[3] = 16'h054D;
assign fc1_node2_c[4] = 16'hF219;
assign fc1_node2_c[5] = 16'h026E;
assign fc1_node2_c[6] = 16'h0D27;
assign fc1_node2_c[7] = 16'h051C;
assign fc1_node2_c[8] = 16'h0B0B;


//FC1_node3
wire signed[15:0] fc1_node3_c[8:0];
assign fc1_node3_c[0] = 16'hEB51;
assign fc1_node3_c[1] = 16'hF29B;
assign fc1_node3_c[2] = 16'hEDD3;
assign fc1_node3_c[3] = 16'h04BA;
assign fc1_node3_c[4] = 16'h0B25;
assign fc1_node3_c[5] = 16'h0383;
assign fc1_node3_c[6] = 16'h04BF;
assign fc1_node3_c[7] = 16'h02D0;
assign fc1_node3_c[8] = 16'h0C5E;


//FC1_node4
wire signed[15:0] fc1_node4_c[8:0];
assign fc1_node4_c[0] = 16'h051C;
assign fc1_node4_c[1] = 16'h0A09;
assign fc1_node4_c[2] = 16'h1748;
assign fc1_node4_c[3] = 16'h0552;
assign fc1_node4_c[4] = 16'h07BA;
assign fc1_node4_c[5] = 16'h0954;
assign fc1_node4_c[6] = 16'h05F8;
assign fc1_node4_c[7] = 16'hF9F7;
assign fc1_node4_c[8] = 16'hF368;


