wire [15:0] FIR_C [99:0];
assign FIR_C[0] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[1] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[2] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[3] = 16'hFFFF;    // -0.00024414062500000000
assign FIR_C[4] = 16'hFFFF;    // -0.00024414062500000000
assign FIR_C[5] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[6] = 16'h0001;    // 0.00024414062500000000
assign FIR_C[7] = 16'h0002;    // 0.00048828125000000000
assign FIR_C[8] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[9] = 16'hFFFF;    // -0.00024414062500000000
assign FIR_C[10] = 16'hFFFC;    // -0.00097656250000000000
assign FIR_C[11] = 16'hFFFD;    // -0.00073242187500000000
assign FIR_C[12] = 16'h0001;    // 0.00024414062500000000
assign FIR_C[13] = 16'h0005;    // 0.00122070312500000000
assign FIR_C[14] = 16'h0006;    // 0.00146484375000000000
assign FIR_C[15] = 16'h0001;    // 0.00024414062500000000
assign FIR_C[16] = 16'hFFFA;    // -0.00146484375000000000
assign FIR_C[17] = 16'hFFF6;    // -0.00244140625000000000
assign FIR_C[18] = 16'hFFFA;    // -0.00146484375000000000
assign FIR_C[19] = 16'h0004;    // 0.00097656250000000000
assign FIR_C[20] = 16'h000E;    // 0.00341796875000000000
assign FIR_C[21] = 16'h000E;    // 0.00341796875000000000
assign FIR_C[22] = 16'h0001;    // 0.00024414062500000000
assign FIR_C[23] = 16'hFFF1;    // -0.00366210937500000000
assign FIR_C[24] = 16'hFFEA;    // -0.00537109375000000000
assign FIR_C[25] = 16'hFFF5;    // -0.00268554687500000000
assign FIR_C[26] = 16'h000C;    // 0.00292968750000000000
assign FIR_C[27] = 16'h001F;    // 0.00756835937500000000
assign FIR_C[28] = 16'h001A;    // 0.00634765625000000000
assign FIR_C[29] = 16'hFFFE;    // -0.00048828125000000000
assign FIR_C[30] = 16'hFFDD;    // -0.00854492187500000000
assign FIR_C[31] = 16'hFFD4;    // -0.01074218750000000000
assign FIR_C[32] = 16'hFFF0;    // -0.00390625000000000000
assign FIR_C[33] = 16'h001F;    // 0.00756835937500000000
assign FIR_C[34] = 16'h003F;    // 0.01538085937500000000
assign FIR_C[35] = 16'h002E;    // 0.01123046875000000000
assign FIR_C[36] = 16'hFFF1;    // -0.00366210937500000000
assign FIR_C[37] = 16'hFFB2;    // -0.01904296875000000000
assign FIR_C[38] = 16'hFFA9;    // -0.02124023437500000000
assign FIR_C[39] = 16'hFFEB;    // -0.00512695312500000000
assign FIR_C[40] = 16'h0051;    // 0.01977539062500000000
assign FIR_C[41] = 16'h008C;    // 0.03417968750000000000
assign FIR_C[42] = 16'h005A;    // 0.02197265625000000000
assign FIR_C[43] = 16'hFFC3;    // -0.01489257812500000000
assign FIR_C[44] = 16'hFF28;    // -0.05273437500000000000
assign FIR_C[45] = 16'hFF15;    // -0.05737304687500000000
assign FIR_C[46] = 16'hFFE8;    // -0.00585937500000000000
assign FIR_C[47] = 16'h0185;    // 0.09497070312500000000
assign FIR_C[48] = 16'h0352;    // 0.20751953125000000000
assign FIR_C[49] = 16'h0481;    // 0.28149414062500000000
assign FIR_C[50] = 16'h0481;    // 0.28149414062500000000
assign FIR_C[51] = 16'h0352;    // 0.20751953125000000000
assign FIR_C[52] = 16'h0185;    // 0.09497070312500000000
assign FIR_C[53] = 16'hFFE8;    // -0.00585937500000000000
assign FIR_C[54] = 16'hFF15;    // -0.05737304687500000000
assign FIR_C[55] = 16'hFF28;    // -0.05273437500000000000
assign FIR_C[56] = 16'hFFC3;    // -0.01489257812500000000
assign FIR_C[57] = 16'h005A;    // 0.02197265625000000000
assign FIR_C[58] = 16'h008C;    // 0.03417968750000000000
assign FIR_C[59] = 16'h0051;    // 0.01977539062500000000
assign FIR_C[60] = 16'hFFEB;    // -0.00512695312500000000
assign FIR_C[61] = 16'hFFA9;    // -0.02124023437500000000
assign FIR_C[62] = 16'hFFB2;    // -0.01904296875000000000
assign FIR_C[63] = 16'hFFF1;    // -0.00366210937500000000
assign FIR_C[64] = 16'h002E;    // 0.01123046875000000000
assign FIR_C[65] = 16'h003F;    // 0.01538085937500000000
assign FIR_C[66] = 16'h001F;    // 0.00756835937500000000
assign FIR_C[67] = 16'hFFF0;    // -0.00390625000000000000
assign FIR_C[68] = 16'hFFD4;    // -0.01074218750000000000
assign FIR_C[69] = 16'hFFDD;    // -0.00854492187500000000
assign FIR_C[70] = 16'hFFFE;    // -0.00048828125000000000
assign FIR_C[71] = 16'h001A;    // 0.00634765625000000000
assign FIR_C[72] = 16'h001F;    // 0.00756835937500000000
assign FIR_C[73] = 16'h000C;    // 0.00292968750000000000
assign FIR_C[74] = 16'hFFF5;    // -0.00268554687500000000
assign FIR_C[75] = 16'hFFEA;    // -0.00537109375000000000
assign FIR_C[76] = 16'hFFF1;    // -0.00366210937500000000
assign FIR_C[77] = 16'h0001;    // 0.00024414062500000000
assign FIR_C[78] = 16'h000E;    // 0.00341796875000000000
assign FIR_C[79] = 16'h000E;    // 0.00341796875000000000
assign FIR_C[80] = 16'h0004;    // 0.00097656250000000000
assign FIR_C[81] = 16'hFFFA;    // -0.00146484375000000000
assign FIR_C[82] = 16'hFFF6;    // -0.00244140625000000000
assign FIR_C[83] = 16'hFFFA;    // -0.00146484375000000000
assign FIR_C[84] = 16'h0001;    // 0.00024414062500000000
assign FIR_C[85] = 16'h0006;    // 0.00146484375000000000
assign FIR_C[86] = 16'h0005;    // 0.00122070312500000000
assign FIR_C[87] = 16'h0001;    // 0.00024414062500000000
assign FIR_C[88] = 16'hFFFD;    // -0.00073242187500000000
assign FIR_C[89] = 16'hFFFC;    // -0.00097656250000000000
assign FIR_C[90] = 16'hFFFF;    // -0.00024414062500000000
assign FIR_C[91] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[92] = 16'h0002;    // 0.00048828125000000000
assign FIR_C[93] = 16'h0001;    // 0.00024414062500000000
assign FIR_C[94] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[95] = 16'hFFFF;    // -0.00024414062500000000
assign FIR_C[96] = 16'hFFFF;    // -0.00024414062500000000
assign FIR_C[97] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[98] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[99] = 16'h0000;    // 0.00000000000000000000
