//conv0 kernel0 coeff
wire signed[15:0] conv0_kernel0_c[4:0];
assign conv0_kernel0_c[0] = 16'hFE51;
assign conv0_kernel0_c[1] = 16'hFDE7;
assign conv0_kernel0_c[2] = 16'hF167;
assign conv0_kernel0_c[3] = 16'hF18A;
assign conv0_kernel0_c[4] = 16'hF561;


//conv0 kernel1 coeff
wire signed[15:0] conv0_kernel1_c[4:0];
assign conv0_kernel1_c[0] = 16'hFCDB;
assign conv0_kernel1_c[1] = 16'hFD2E;
assign conv0_kernel1_c[2] = 16'h0548;
assign conv0_kernel1_c[3] = 16'h007E;
assign conv0_kernel1_c[4] = 16'h03A1;


//conv0 kernel2 coeff
wire signed[15:0] conv0_kernel2_c[4:0];
assign conv0_kernel2_c[0] = 16'hF7B1;
assign conv0_kernel2_c[1] = 16'hF5C7;
assign conv0_kernel2_c[2] = 16'hEF4F;
assign conv0_kernel2_c[3] = 16'hF27A;
assign conv0_kernel2_c[4] = 16'hF6C4;


//conv0 kernel3 coeff
wire signed[15:0] conv0_kernel3_c[4:0];
assign conv0_kernel3_c[0] = 16'h00E6;
assign conv0_kernel3_c[1] = 16'h0221;
assign conv0_kernel3_c[2] = 16'h02E5;
assign conv0_kernel3_c[3] = 16'hF9AC;
assign conv0_kernel3_c[4] = 16'hFBBE;


//conv0 kernel4 coeff
wire signed[15:0] conv0_kernel4_c[4:0];
assign conv0_kernel4_c[0] = 16'h0E79;
assign conv0_kernel4_c[1] = 16'h1837;
assign conv0_kernel4_c[2] = 16'h1113;
assign conv0_kernel4_c[3] = 16'h14A7;
assign conv0_kernel4_c[4] = 16'h0A74;


//conv1 kernel0_0 coeff
wire signed[15:0] conv1_kernel0_0_c[4:0];
assign conv1_kernel0_0_c[0] = 16'h0706;
assign conv1_kernel0_0_c[1] = 16'h1182;
assign conv1_kernel0_0_c[2] = 16'h0CAF;
assign conv1_kernel0_0_c[3] = 16'h0733;
assign conv1_kernel0_0_c[4] = 16'hFF9A;


//conv1 kernel0_1 coeff
wire signed[15:0] conv1_kernel0_1_c[4:0];
assign conv1_kernel0_1_c[0] = 16'hFD8F;
assign conv1_kernel0_1_c[1] = 16'h01C5;
assign conv1_kernel0_1_c[2] = 16'hFD16;
assign conv1_kernel0_1_c[3] = 16'hFE06;
assign conv1_kernel0_1_c[4] = 16'hFD49;


//conv1 kernel0_2 coeff
wire signed[15:0] conv1_kernel0_2_c[4:0];
assign conv1_kernel0_2_c[0] = 16'h039A;
assign conv1_kernel0_2_c[1] = 16'h0F87;
assign conv1_kernel0_2_c[2] = 16'h16AD;
assign conv1_kernel0_2_c[3] = 16'h0D15;
assign conv1_kernel0_2_c[4] = 16'h02B3;


//conv1 kernel0_3 coeff
wire signed[15:0] conv1_kernel0_3_c[4:0];
assign conv1_kernel0_3_c[0] = 16'h01DF;
assign conv1_kernel0_3_c[1] = 16'h010F;
assign conv1_kernel0_3_c[2] = 16'h0257;
assign conv1_kernel0_3_c[3] = 16'hFDA1;
assign conv1_kernel0_3_c[4] = 16'hFDE6;


//conv1 kernel0_4 coeff
wire signed[15:0] conv1_kernel0_4_c[4:0];
assign conv1_kernel0_4_c[0] = 16'hFDB2;
assign conv1_kernel0_4_c[1] = 16'hFBE9;
assign conv1_kernel0_4_c[2] = 16'hFB4B;
assign conv1_kernel0_4_c[3] = 16'hFE40;
assign conv1_kernel0_4_c[4] = 16'hFEB8;


//conv1 kernel1_0 coeff
wire signed[15:0] conv1_kernel1_0_c[4:0];
assign conv1_kernel1_0_c[0] = 16'h04A3;
assign conv1_kernel1_0_c[1] = 16'h03D4;
assign conv1_kernel1_0_c[2] = 16'h0442;
assign conv1_kernel1_0_c[3] = 16'hFFBB;
assign conv1_kernel1_0_c[4] = 16'hFED0;


//conv1 kernel1_1 coeff
wire signed[15:0] conv1_kernel1_1_c[4:0];
assign conv1_kernel1_1_c[0] = 16'h0109;
assign conv1_kernel1_1_c[1] = 16'h04E5;
assign conv1_kernel1_1_c[2] = 16'h01E5;
assign conv1_kernel1_1_c[3] = 16'h006D;
assign conv1_kernel1_1_c[4] = 16'h031D;


//conv1 kernel1_2 coeff
wire signed[15:0] conv1_kernel1_2_c[4:0];
assign conv1_kernel1_2_c[0] = 16'h0495;
assign conv1_kernel1_2_c[1] = 16'hFFFF;
assign conv1_kernel1_2_c[2] = 16'h0373;
assign conv1_kernel1_2_c[3] = 16'h00B2;
assign conv1_kernel1_2_c[4] = 16'h0131;


//conv1 kernel1_3 coeff
wire signed[15:0] conv1_kernel1_3_c[4:0];
assign conv1_kernel1_3_c[0] = 16'h007E;
assign conv1_kernel1_3_c[1] = 16'h0224;
assign conv1_kernel1_3_c[2] = 16'h01B6;
assign conv1_kernel1_3_c[3] = 16'h029D;
assign conv1_kernel1_3_c[4] = 16'h018F;


//conv1 kernel1_4 coeff
wire signed[15:0] conv1_kernel1_4_c[4:0];
assign conv1_kernel1_4_c[0] = 16'hD72B;
assign conv1_kernel1_4_c[1] = 16'h0E22;
assign conv1_kernel1_4_c[2] = 16'h138F;
assign conv1_kernel1_4_c[3] = 16'h12B8;
assign conv1_kernel1_4_c[4] = 16'h0C69;


